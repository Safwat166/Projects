package pack ;
    import uvm_pkg::* ;
    `include "uvm_macros.svh"
    `include "classes/sequence_item.sv"
    `include "classes/sequence.sv"
    `include "classes/sequencer.sv"
    `include "classes/driver.sv"
    `include "classes/monitor.sv"
    `include "classes/agent.sv"
    `include "classes/scoreboard.sv"
    `include "classes/enviroment.sv"
    `include "classes/test.sv"
endpackage : pack