package pack ;
    import uvm_pkg::* ;
    `include    "uvm_macros.svh"
    `include    "Classes/Sequence_Item_Class.sv"
    `include    "Classes/Sequence_Class.sv"
    `include    "Classes/Driver_Class.sv"
    `include    "Classes/Monitor_Class.sv"
    `include    "Classes/Sequencer_Class.sv"
    `include    "Classes/Agent_Class.sv"
    `include    "Classes/Scoreboard_Class.sv"
    `include    "Classes/Env_Class.sv"
    `include    "Classes/Test_Class.sv"
endpackage : pack