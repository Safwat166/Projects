package pack ;
    `include    "Classes/Transaction_Class.sv"
    `include    "Classes/Driver_Class.sv"
    `include    "Classes/Monitor_Class.sv"
    `include    "Classes/Scoreboard_Class.sv"
    `include    "Classes/Sequencer_Class.sv"
    `include    "Classes/Env_Class.sv"
endpackage